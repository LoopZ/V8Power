vline [flaggor]

Ritar en linje.

    [inga]      Ritar en lokal, enkel dum linje p� aktuell rad.
    /K n        Anv�nd n ist�llet f�r ramtecken f�r att identifiera ramar.
    single      Ritar en enkel linje.
    double      Ritar en dubbel linje.
    hidden      Ritar en osynlig dum linje.
    dumb        Ritar en dum linje utan h�nsyn taget till vad som redan finns.

    tba         (Fortfarande under utveckling, mer kommer att annonseras)

