vmode [flaggor]

S�tt och fr�ga efter aktuellt textl�ge.

    [inga]      Skriver ut aktuellt videol�ge och typsnitt till STDOUT.
    VESA        Skriver ut en lista �ver VESA-l�gen till STDOUT.
    l�ge        S�tt aktuellt videol�ge. (0-0xffff) eller l�gesetikett
                med valfri typsnittsinst�llning

                L�gen:  BW40    Svart/vitt 40 kolumner (ocks� B40).
                        BW80    Svart/vitt 80 kolumner (ocks� B80, BW).
                        CO40    F�rg 40 kolumner (ocks� C40).
                        CO80    F�rg 80 kolumner (ocks� C80, COLOR).
                        MONO    Monokrom 80 kolumner.

                Typsnitt:  Font8   V�ljer 8x8 ROM-typsnitt. (ocks� F8)
                           Font14  V�ljer 8x14 EGA ROM-typsnitt. (ocks� F14)
                           Font16  V�ljer 8x16 VGA ROM-typsnitt. (ocks� F16)

