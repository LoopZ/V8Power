vcls [flaggor]

Rensa sk�rmen, omr�det eller rad.

    [inga]      Rensa sk�rmen med aktuellt textattribut.
    n           S�tt textattribut till n.
    /A n        S�tt textattribut till n.
    /B f�rg     S�tt textattribut f�r bakgrunden till f�rg (eller v�rde).
    /F f�rg     S�tt textattribut f�r f�rgrunden till f�rg (eller v�rde).
    /G          Globak sk�rmrensning. (Standard)
    /L          Lokal sk�rmrensning. Detekterar dess omgivningar och rensar
                endast den. Troligtvis en ruta eller rad eller n�got. Du m�ste
		inte anv�nda denna flagga d� du helt enkelt kan rita om rutan.
    /K n        Anv�nd n ist�llet f�r ramtecken f�r att identifiera ramar.
    TEXT        Rensar endast texten. L�mna alla f�rger intakta och hoppa �ver
                deras f�rgattribut.
    EOL         Rensar endast fr�n mark�ren till slutet p� raden.
    /C kod      Rensa genom att fylla med ASCII-teckenkod.
    /X kolumn   Absolut sk�rmkolumn att b�rja rensa p�.
    /Y rad      Absolut sk�rmrad att b�rja resan p�
    /W bredd    Total bredd p� omr�de att rensa.
    /H h�jd     Total h�jd p� omr�de att rensa.
