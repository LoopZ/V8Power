vask [flaggor]

Fr�ga efter textinmatning.

    [inga]      Anv�nd identifierade inst�llningar f�r inmatning.
    [text]      F�rinst�ll redigerad text.
    /A n        S�tt textattribut till n.
    /B f�rg     S�tt textattribut f�r bakgrund till f�rg (eller v�rde).
    /F f�rg     S�tt textattribut f�r f�rgrund till f�rg (eller v�rde).
    /G          Mata in text globalt och ignorera alla ramar.
    /L          Mata in text lokalt med h�nsyn tagen till ramar. (STANDARD)
    /K n        Anv�nd n ist�llet f�r ramtecken f�r att identifiera ramar.
    /C          N�r angivet och Ctrl-C trycks, avsluta med
                errorlevel 200 och returnera standardv�rdet.
    /W bredd    �sidos�tt standardbredd f�r raden.
                (standard �r fr�n mark�ren till slutet p� raden)
    /T fil ID   Sl� upp ID i fil och behandla den som en kommandoradsparameter.
                Ytterligare parametrar som f�ljer p� denna flagga anv�nds f�r
		att populera variablerna %1-%9 i textstr�ngen.
    /D sekunder F�rdr�jning i sekunder att v�nta innan tidsgr�nsen f�r
                inmatningsf�rfr�gan l�per ut och returnera det inledande
		standardv�rdet. (returnerar errorlevel 1)

    tba         (Fortfarande under utveckling, mer kommer att annonseras)

