vgotoxy [flaggor]

Flytta eller fr�ga efter mark�rposition.

    [inga]      Utf�r ingen �tg�rd
    /Q x        Fr�ga om aktuell X eller Y position f�r mark�ren och matar
    /Q y        ut den till STDOUT.
    /X kolumn   Flytta mark�r till kolumn.
    /Y rad      Flytta mark�r till rad.
    /G          Flytta mark�r baserat p� hela sk�rmen. (standard)
    /L          Flytta mark�r baserat p� dess omgivning.
    /K n        Anv�nd n ist�llet f�r ramtecken f�r att identifierar ramar.
    direction   Flytta mark�r upp, ner, v�nster eller h�ger ett steg.
    shift       Flytta mark�r till f�reg�ende eller n�sta position och �ndra
                rader om det beh�vs.
    position    Flytta mark�r till
                    SOP (B�rjan av sidan),
                    EOP (Slutet av sidan),
                    SOR (B�rjan av raden),
                    EOR (Slutet av raden),
                    SOL (B�rjan av text p� rad),
                    EOL (Slutet av text p� rad),
                    SOT (B�rjan av all text) eller
                    EOT (Slutet av all text).
