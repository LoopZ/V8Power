vcursor [flaggor]

�ndra eller fr�ga om mark�rstorlek och form.

    [inga]      Skriver ut aktuell mark�rform till STDOUT.
    n           S�tter aktuell mark�rform till n.
    HIDE        G�mmer mark�ren.
    SMALL       S�tter en liten mark�r.
    HALF        S�tter mark�ren till halv texth�jden.
    FULL        S�tter mark�ren till hela texth�jden.

Notera: �ven om detta verktyg �r fullt kompatibelt med DOSBox finns det
inget s�tt att lagra aktuell mark�rform. Se exemplen f�r hur du kringg�r
detta problem. Detta verktyg har hellet inte n�gon effekt i en
Windows-terminal.
