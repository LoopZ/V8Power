vdelay [ms]

Enkel f�rdr�jning i millisekunder.

    [inga]      Standard f�rdr�jning �r 1000ms (1 sekund).
    ms          F�rdr�jning i ms millisekunder. (0-65535, 0x0000-0xffff)
    /D          Identifiera f�rdr�jningsmetod. (Inte kompatibelt med VirtualBox)
    /S          Anv�nd s�ker timer f�r allm�nt bruk. (Standard)
    /I          Anv�nd h�gprecisions timeravbrott. (Inte kompatibelt med
                VirtualBox)
