vfont [flaggor]
L�s tillf�lligt in ett bitmapstypsnitt f�r textl�ge.

    fil         L�s in typsnittsfil.
    /F n fil    Om aktuellt typsnitt har n (nummer, EGA eller VGA) rader
                l�s d� in typsnittsfilen. Kan kedjas f�r olika uppl�sningar.
    /D          L�s in standardtypsnitt f�r aktuell uppl�sning.

   tba         (Fortfarande under utveckling, mer kommer att annonseras)

