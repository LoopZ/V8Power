verrlvl [flaggor]

S�tt aktuell errorlevel. Mestadels f�r att testa logiken i kommandofiler.

    [inga]      S�tter errorlevel till 0
    n           S�tter errorlevel till n (0-255)

