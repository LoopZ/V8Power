vprogres [flaggor]

Rita en f�rloppsindikator p� aktuell position utan att flytta mark�ren.

    [inga]      Rita en f�rloppsindikator med 0%.
    /A n        S�tt textattribut till n.
    /B f�rg     S�tt textattribut f�r bakgrunden till f�rg (eller v�rde).
    /F f�rg     S�tt textattribut f�r f�rgrunden till f�rg (eller v�rde).
    /W bredd    �sidos�tt standard bredd f�r f�rloppindikatorn.
                (standard �r fr�n mark�ren till radslutet)
    /K n        Anv�nd n ist�llet f�r ramtecken f�r att identifiera ramar.
    v�rde       S�tter v�rdet i procent f�r f�rloppet.
    off         Visa inte procentantal.
    justering   Procentnummer till v�nster, centrerat (Standard) eller till
                h�ger om f�rloppsindikatorn.
    OF max      Ber�kna procentandel av max. Till exempel 5 av 7.

