vframe [flaggor]

Rita en f�nsterruta och flytta in mark�ren till dess �vre v�nstra h�rn.

    [inga]      Rita en ruta som t�cker hela sk�rmen.
    /A n        S�tt textattribut till n.
    /B f�rg     S�tt textattribut f�r bakgrunden till f�rg (eller v�rde).
    /F f�rg     S�tt textattribut f�r f�rgrunden till f�rg (eller v�rde).
    /X kolumn   B�rja rutan p� sk�rmkolumn kolumn.
    /Y rad      B�rja rutan p� sk�rmrad rad.
    /W bredd    Total bredd f�r rutan.
    /H h�jd     Total h�jd f�r rutan.
    /C          Centrerar rutan horisontellt och vertikalt.
    /T fil ID   Sl� upp ID i fil och behandla det som en kommandoradsparameter.
                Resterande parametrar som f�ljer denna flagga anv�nds f�r att
		populera variablerna %1-%9 i textstr�ngen.
    /P n        S�tter ett osynligt utfyllnadstecken n f�r textrutor och
                alternativrutor.
    style       Boxstilar �r Single, Double, SingleSides, DoubleSides
                och Hidden.
    shadow      L�gg till en 3D-skugga.
    textbox     Rita en ram i textboxstil med lite utfyllnad och marginaler.
    optionbox   Rita en alternativbox i g�md stil f�r alternativ inuti en ram.
